module registerfile(
    
);
    
endmodule //registerfile