module mem_ctrl (
    input   wire    clk,
    input   wire    rst,
    input   wire    rdy,
    
    input   wire    rollback, // 1 means Reorder Buffer need rollback

    input   wire    [7:0]   data_in, // for write
    output  


);
    
endmodule //mem_ctrl
