module mem_ctrl (
    input   wire    clk,
    input   wire    rst,
    input   wire    rdy,
    
);
    
endmodule //mem_ctrl
